module fetch();

endmodule

