module decode();


endmodule

