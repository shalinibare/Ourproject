module cpu_mem();

endmodule

