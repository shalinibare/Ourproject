module imm_extender_tb()


endmodule
