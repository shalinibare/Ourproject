module Branch_calc_tb();


endmodule
