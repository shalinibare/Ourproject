module Forwarding_Unit();

endmodule

