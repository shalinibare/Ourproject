//Module to initiate DMA controller transactions (Read layer inputs, images,
//etc.)
module DMA_FSM();


endmodule

