module cpu_top();


endmodule

