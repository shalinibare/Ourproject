module Register_File_tb();


endmodule

