module Control_tb();


endmodule

