module execute();


endmodule

