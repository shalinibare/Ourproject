module memory_controller_tb ();
    localparam  DATA_WIDTH=32;
    localparam  ADDR_WIDTH=16;
    localparam  TEST_CASE=100;
    
endmodule